netcdf TestData {
dimensions:
    x = 10 ;
    y = 10 ;
    time = 4 ;
variables:
    int x(x) ;
    int y(y) ;
    float z(x, y) ;
    float h(time, y, x) ;
    float hu(time, y, x) ;
    float hv(time, y, x) ;
    float b(y, x) ;
data:
   x = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9 ;
   y = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9 ;
   z = 
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
   b = 
        10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
        20, 20, 20, 20, 20, 20, 20, 20, 20, 20,
        30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
        40, 40, 40, 40, 40, 40, 40, 40, 40, 40,
        50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
        60, 60, 60, 60, 60, 60, 60, 60, 60, 60,
        70, 70, 70, 70, 70, 70, 70, 70, 70, 70,
        80, 80, 80, 80, 80, 80, 80, 80, 80, 80,
        90, 90, 90, 90, 90, 90, 90, 90, 90, 90,
        100, 100, 100, 100, 100, 100, 100, 100, 100, 100 ;
        
}
